`include "CPU\\InstructionDecoder\\InstructionDecoder.v"
`timescale 100ns/100ns

module tb;
    reg [15:0] Instruction;

    wire [15:0] FS, BranchOffset;
    wire [3:0] srcA, dstA;
    wire [1:0] As;
    wire Ad, BW, OneOp;

    InstructionDecoder uut(
        .Instruction(Instruction),
        .FS(FS), .BranchOffset(BranchOffset),
        .srcA(srcA), .dstA(dstA),
        .As(As), .Ad(Ad), .BW(BW), .OneOp(OneOp)
    );

    initial begin
        $dumpfile("InstructionDecoder.vcd");
        $dumpvars(0, tb);
        // Dump Instructions Here
        Instruction = 16'h1004; #10;
        Instruction = 16'h1025; #10;
        Instruction = 16'h1036; #10;
        Instruction = 16'h1017; #10;
        Instruction = 16'h1044; #10;
        Instruction = 16'h1065; #10;
        Instruction = 16'h1076; #10;
        Instruction = 16'h1057; #10;
        Instruction = 16'h1088; #10;
        Instruction = 16'h10A9; #10;
        Instruction = 16'h10BA; #10;
        Instruction = 16'h109B; #10;
        Instruction = 16'h110C; #10;
        Instruction = 16'h112D; #10;
        Instruction = 16'h113E; #10;
        Instruction = 16'h111F; #10;
        Instruction = 16'h114C; #10;
        Instruction = 16'h116D; #10;
        Instruction = 16'h117E; #10;
        Instruction = 16'h115F; #10;
        Instruction = 16'h1184; #10;
        Instruction = 16'h11A6; #10;
        Instruction = 16'h11B8; #10;
        Instruction = 16'h1198; #10;
        Instruction = 16'h1205; #10;
        Instruction = 16'h1226; #10;
        Instruction = 16'h1237; #10;
        Instruction = 16'h1230; #10;
        Instruction = 16'h121B; #10;
        Instruction = 16'h1245; #10;
        Instruction = 16'h1266; #10;
        Instruction = 16'h1277; #10;
        Instruction = 16'h1270; #10;
        Instruction = 16'h125B; #10;
        Instruction = 16'h1284; #10;
        Instruction = 16'h12A5; #10;
        Instruction = 16'h12B6; #10;
        Instruction = 16'h12B0; #10;
        Instruction = 16'h1297; #10;
        Instruction = 16'h1300; #10;
        Instruction = 16'h2009; #10;
        Instruction = 16'h2008; #10;
        Instruction = 16'h2407; #10;
        Instruction = 16'h2406; #10;
        Instruction = 16'h2805; #10;
        Instruction = 16'h2C04; #10;
        Instruction = 16'h33F9; #10;
        Instruction = 16'h37F8; #10;
        Instruction = 16'h3BF7; #10;
        Instruction = 16'h3FF6; #10;
        Instruction = 16'h4407; #10;
        Instruction = 16'h4588; #10;
        Instruction = 16'h4629; #10;
        Instruction = 16'h47AA; #10;
        Instruction = 16'h483B; #10;
        Instruction = 16'h49BC; #10;
        Instruction = 16'h403D; #10;
        Instruction = 16'h4A1E; #10;
        Instruction = 16'h4B9F; #10;
        Instruction = 16'h4845; #10;
        Instruction = 16'h49C6; #10;
        Instruction = 16'h4A67; #10;
        Instruction = 16'h4BE8; #10;
        Instruction = 16'h4C79; #10;
        Instruction = 16'h4DFA; #10;
        Instruction = 16'h407B; #10;
        Instruction = 16'h4E5C; #10;
        Instruction = 16'h4FDD; #10;
        Instruction = 16'h5407; #10;
        Instruction = 16'h5588; #10;
        Instruction = 16'h5629; #10;
        Instruction = 16'h57AA; #10;
        Instruction = 16'h583B; #10;
        Instruction = 16'h59BC; #10;
        Instruction = 16'h503D; #10;
        Instruction = 16'h5A1E; #10;
        Instruction = 16'h5B9F; #10;
        Instruction = 16'h5845; #10;
        Instruction = 16'h59C6; #10;
        Instruction = 16'h5A67; #10;
        Instruction = 16'h5BE8; #10;
        Instruction = 16'h5C79; #10;
        Instruction = 16'h5DFA; #10;
        Instruction = 16'h507B; #10;
        Instruction = 16'h5E5C; #10;
        Instruction = 16'h5FDD; #10;
        Instruction = 16'h6407; #10;
        Instruction = 16'h6588; #10;
        Instruction = 16'h6629; #10;
        Instruction = 16'h67AA; #10;
        Instruction = 16'h683B; #10;
        Instruction = 16'h69BC; #10;
        Instruction = 16'h603D; #10;
        Instruction = 16'h6A1E; #10;
        Instruction = 16'h6B9F; #10;
        Instruction = 16'h6845; #10;
        Instruction = 16'h69C6; #10;
        Instruction = 16'h6A67; #10;
        Instruction = 16'h6BE8; #10;
        Instruction = 16'h6C79; #10;
        Instruction = 16'h6DFA; #10;
        Instruction = 16'h607B; #10;
        Instruction = 16'h6E5C; #10;
        Instruction = 16'h6FDD; #10;
        Instruction = 16'h7407; #10;
        Instruction = 16'h7588; #10;
        Instruction = 16'h7629; #10;
        Instruction = 16'h77AA; #10;
        Instruction = 16'h783B; #10;
        Instruction = 16'h79BC; #10;
        Instruction = 16'h703D; #10;
        Instruction = 16'h7A1E; #10;
        Instruction = 16'h7B9F; #10;
        Instruction = 16'h7845; #10;
        Instruction = 16'h79C6; #10;
        Instruction = 16'h7A67; #10;
        Instruction = 16'h7BE8; #10;
        Instruction = 16'h7C79; #10;
        Instruction = 16'h7DFA; #10;
        Instruction = 16'h707B; #10;
        Instruction = 16'h7E5C; #10;
        Instruction = 16'h7FDD; #10;
        Instruction = 16'h8407; #10;
        Instruction = 16'h8588; #10;
        Instruction = 16'h8629; #10;
        Instruction = 16'h87AA; #10;
        Instruction = 16'h883B; #10;
        Instruction = 16'h89BC; #10;
        Instruction = 16'h803D; #10;
        Instruction = 16'h8A1E; #10;
        Instruction = 16'h8B9F; #10;
        Instruction = 16'h8845; #10;
        Instruction = 16'h89C6; #10;
        Instruction = 16'h8A67; #10;
        Instruction = 16'h8BE8; #10;
        Instruction = 16'h8C79; #10;
        Instruction = 16'h8DFA; #10;
        Instruction = 16'h807B; #10;
        Instruction = 16'h8E5C; #10;
        Instruction = 16'h8FDD; #10;
        Instruction = 16'h9407; #10;
        Instruction = 16'h9588; #10;
        Instruction = 16'h9629; #10;
        Instruction = 16'h97AA; #10;
        Instruction = 16'h983B; #10;
        Instruction = 16'h99BC; #10;
        Instruction = 16'h903D; #10;
        Instruction = 16'h9A1E; #10;
        Instruction = 16'h9B9F; #10;
        Instruction = 16'h9845; #10;
        Instruction = 16'h99C6; #10;
        Instruction = 16'h9A67; #10;
        Instruction = 16'h9BE8; #10;
        Instruction = 16'h9C79; #10;
        Instruction = 16'h9DFA; #10;
        Instruction = 16'h907B; #10;
        Instruction = 16'h9E5C; #10;
        Instruction = 16'h9FDD; #10;
        Instruction = 16'hA407; #10;
        Instruction = 16'hA588; #10;
        Instruction = 16'hA629; #10;
        Instruction = 16'hA7AA; #10;
        Instruction = 16'hA83B; #10;
        Instruction = 16'hA9BC; #10;
        Instruction = 16'hA03D; #10;
        Instruction = 16'hAA1E; #10;
        Instruction = 16'hAB9F; #10;
        Instruction = 16'hA845; #10;
        Instruction = 16'hA9C6; #10;
        Instruction = 16'hAA67; #10;
        Instruction = 16'hABE8; #10;
        Instruction = 16'hAC79; #10;
        Instruction = 16'hADFA; #10;
        Instruction = 16'hA07B; #10;
        Instruction = 16'hAE5C; #10;
        Instruction = 16'hAFDD; #10;
        Instruction = 16'hB407; #10;
        Instruction = 16'hB588; #10;
        Instruction = 16'hB629; #10;
        Instruction = 16'hB7AA; #10;
        Instruction = 16'hB83B; #10;
        Instruction = 16'hB9BC; #10;
        Instruction = 16'hB03D; #10;
        Instruction = 16'hBA1E; #10;
        Instruction = 16'hBB9F; #10;
        Instruction = 16'hB845; #10;
        Instruction = 16'hB9C6; #10;
        Instruction = 16'hBA67; #10;
        Instruction = 16'hBBE8; #10;
        Instruction = 16'hBC79; #10;
        Instruction = 16'hBDFA; #10;
        Instruction = 16'hB07B; #10;
        Instruction = 16'hBE5C; #10;
        Instruction = 16'hBFDD; #10;
        Instruction = 16'hC407; #10;
        Instruction = 16'hC588; #10;
        Instruction = 16'hC629; #10;
        Instruction = 16'hC7AA; #10;
        Instruction = 16'hC83B; #10;
        Instruction = 16'hC9BC; #10;
        Instruction = 16'hC03D; #10;
        Instruction = 16'hCA1E; #10;
        Instruction = 16'hCB9F; #10;
        Instruction = 16'hC845; #10;
        Instruction = 16'hC9C6; #10;
        Instruction = 16'hCA67; #10;
        Instruction = 16'hCBE8; #10;
        Instruction = 16'hCC79; #10;
        Instruction = 16'hCDFA; #10;
        Instruction = 16'hC07B; #10;
        Instruction = 16'hCE5C; #10;
        Instruction = 16'hCFDD; #10;
        Instruction = 16'hD407; #10;
        Instruction = 16'hD588; #10;
        Instruction = 16'hD629; #10;
        Instruction = 16'hD7AA; #10;
        Instruction = 16'hD83B; #10;
        Instruction = 16'hD9BC; #10;
        Instruction = 16'hD03D; #10;
        Instruction = 16'hDA1E; #10;
        Instruction = 16'hDB9F; #10;
        Instruction = 16'hD845; #10;
        Instruction = 16'hD9C6; #10;
        Instruction = 16'hDA67; #10;
        Instruction = 16'hDBE8; #10;
        Instruction = 16'hDC79; #10;
        Instruction = 16'hDDFA; #10;
        Instruction = 16'hD07B; #10;
        Instruction = 16'hDE5C; #10;
        Instruction = 16'hDFDD; #10;
        Instruction = 16'hE407; #10;
        Instruction = 16'hE588; #10;
        Instruction = 16'hE629; #10;
        Instruction = 16'hE7AA; #10;
        Instruction = 16'hE83B; #10;
        Instruction = 16'hE9BC; #10;
        Instruction = 16'hE03D; #10;
        Instruction = 16'hEA1E; #10;
        Instruction = 16'hEB9F; #10;
        Instruction = 16'hE845; #10;
        Instruction = 16'hE9C6; #10;
        Instruction = 16'hEA67; #10;
        Instruction = 16'hEBE8; #10;
        Instruction = 16'hEC79; #10;
        Instruction = 16'hEDFA; #10;
        Instruction = 16'hE07B; #10;
        Instruction = 16'hEE5C; #10;
        Instruction = 16'hEFDD; #10;
        Instruction = 16'hF407; #10;
        Instruction = 16'hF588; #10;
        Instruction = 16'hF629; #10;
        Instruction = 16'hF7AA; #10;
        Instruction = 16'hF83B; #10;
        Instruction = 16'hF9BC; #10;
        Instruction = 16'hF03D; #10;
        Instruction = 16'hFA1E; #10;
        Instruction = 16'hFB9F; #10;
        Instruction = 16'hF845; #10;
        Instruction = 16'hF9C6; #10;
        Instruction = 16'hFA67; #10;
        Instruction = 16'hFBE8; #10;
        Instruction = 16'hFC79; #10;
        Instruction = 16'hFDFA; #10;
        Instruction = 16'hF07B; #10;
        Instruction = 16'hFE5C; #10;
        Instruction = 16'hFFDD; #10;
        $finish;
    end
endmodule